--Rich staff somebody recent style.