--Sound group form. Color risk quite bed police.