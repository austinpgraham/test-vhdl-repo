--Message education message money.