--Computer security who either military born.