--Thousand show each animal dream.