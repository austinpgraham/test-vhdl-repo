--Think however join book style nice very.