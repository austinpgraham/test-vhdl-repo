--Less song measure sell.