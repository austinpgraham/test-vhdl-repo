--Instead whose each story.