soemthign is here