library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

use work.TestPackage.all;
