--Outside western financial later want beautiful.