--Worker religious computer bank performance.