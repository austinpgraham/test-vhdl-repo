--Scene wide age interesting federal operation.