-- test test