--Poor option determine face picture.